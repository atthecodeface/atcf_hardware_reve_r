/** @copyright (C) 2016-2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_csrs_minimal.cdl
 * @brief  Control/status registers for a minimal RISC-V implementation
 *
 * This file contains a module that implements the in-CPU CSRs
 * required by a RISC-V implementation.
 */

/*a Includes */
include "reve_r_internal_types.h"

/*a Types */
/*t t_csr_write */
typedef struct {
    bit     enable      "Asserted if a CSR write is in progress";
    bit[32] data_mask   "Bits to keep";
    bit[32] data_set    "Bits to set";
} t_csr_write;

/*t t_csr_combs */
typedef struct {
    bit[32] ustatus;
    bit[32] utvec;
    bit[32] uip;
    bit[32] uie;

    bit[32] mstatus;
    bit[32] mtvec;
    bit[32] mip;
    bit[32] mie;

    bit[32] dcsr;
} t_csr_combs;

/*t t_mode_combs */
typedef struct {
    bit d;
    bit m;
    bit s;
    bit u;
} t_mode_combs;

/*a Module */
module reve_r_csrs( clock clk                                   "Free-running clock",
                     clock riscv_clk                             "Clk gated by riscv_clk_enable - provide for single clock gate outside the module",
                     input bit riscv_clk_enable                  "RISC-V clock enable",
                     input bit reset_n                           "Active low reset",
                     input t_riscv_irqs          irqs            "Interrupts in to the CPU",
                     input t_riscv_csr_access    csr_access      "RISC-V CSR access, combinatorially decoded",
                     output t_riscv_csr_data     csr_data        "CSR respone (including read data), from the current @a csr_access",
                     input t_riscv_csr_controls  csr_controls    "Control signals to update the CSRs",
                     output t_riscv_csrs         csrs            "CSR values"
    )
"""
This module implements a minimal set of RISC-V CSRs, as per v2.1 (May
2016) of the RISC-V instruction set manual user level ISA and v1.9.1
of the privilege architecture (Nov 2016), with the exception that
MTIME has been removed (as this seems to be the correct thing to do).

The privilege specifcation (v1.10) indicates:

* meip is read-only and is derived from the external irq in to this module

* mtip is read-only, cleared by writing to the memory-mapped timer comparator

* msip is read-write in a memory-mapped register somewhere

Hence the irqs structure must provide these three signals


Minimal CSRs as only machine mode and debug mode are supported.
In debug mode every register access is supported.
In machine mode then every register EXCEPT access to ??? is supported.

Given machine mode is the only mode supported:

* there are no SEI and UEI interrupt pins in to this module

* SEIP and UEIP are not supported

* STIP and UTIP are not supported

* SSIP and USIP are not supported

* mstatus.SIE and mstatus.UIE (and previous versions) are hardwired to 0

* mstatus.SPP and mstatus.UPP are hardwired to 0

The mip (machine interrupt pending register) therefore is:

{20b0, MEIP, 3b0, MTIP, 3b0, MSIP, 3b0}

The mie (machine interrupt enable register) is:

{20b0, MEIE, 3b0, MTIE, 3b0, MSIE, 3b0}


The instruction to the pipeline to request an interrupt (which is only
taken if an instruction is in uncommitted in the execution stage) must be generated using the
execution mode and the interrupt enable bits and the interrupt pending
bits.

Hence the 'take interrupt' is (mip & mie) != 0 && mstatus.MIE && (current mode >= machine mode) && (current mode != debug mode).

The required priority order is:

external interrupts, software interrupts, timer interrupts

If an instruction has been committed then it may trap, and the trap
will occur prior to an interrupt which happens after the commit
point. In this case there will be a trap, and the trapped instruction
will be fetched, and then an interrupt can be taken.

When an interrupt is taken the following occurs:

* MPP <= current execution mode (must be machine mode, as debug mode is not interruptible)

* mstatus.MPIE <= mstatus.MIE

Note that WFI should wait independent of mstatus.MIE for (mip & mie) != 0 (given machine mode only)
In debug mode WFI should be a NOP.

WFI may always be a NOP.


User mode interrupts
--------------------

For user mode interrupts there has to be support for delegating an interrupt to user mode - hence the medeleg and mideleg need support (read/write)

User mode interrupts are disabled if mstatus.uie is clear

When an interrupt/exception is delegated to user mode uepc/ucause/utval/mstatus.upie are set to the address, cause etc and mstatus.uie at the interrupt/exception
mstatus.uie is a bit of mstatus that is CLEARED on a user interrupt/exception, and which is set to mstatus.upie on uret; mstatus.upie is then set

uscratch is a 32-bit register for use in the trap handler (and outside it too, if necessary)

utvec is a user vector base for vectored user interrupts

mstatus.uie and mstatus.upie are visible (and only these 2 bits) in 'ustatus'

On uret, uepc/ucause/utval can be cleared (i.e. they are guaranteed to be invalid outside of a user trap handler). mstatus.uie become mstatus.upie; mstatus.upie is set; pc becomes mstatus.uepc

The following CSRs should therefore be supplied for user mode interrupts: ustatus, uie, utvec, uscratch, uepc, ucause, utval, uip.
"""
{

    /*b State and combs
     */
    default clock clk;
    default reset active_low reset_n;
    clocked bit keep_clk = 0 "State bit to ensure that 'clk' is kept - can be used be other versions for state updates etc";
    default clock riscv_clk;
    clocked t_riscv_csrs csrs={*=0};
    comb t_csr_combs  csr_combs;
    comb t_csr_write  csr_write;
    comb t_mode_combs ret_combs  "Breakout for xRET";
    comb t_mode_combs trap_combs "Breakout for valid trap to mode";

    /*b Clock 'clk' state
     */
    clk_state :{
        keep_clk <= 0;
    }

    /*b CSR comb bundling
     */
    csr_bundling """
    """: {
        csr_combs.mstatus = bundle(csrs.mstatus.sd,
                         8b0,
                         csrs.mstatus.tsr,
                         csrs.mstatus.tw,
                         csrs.mstatus.tvm,
                         csrs.mstatus.mxr,
                         csrs.mstatus.sum,
                         csrs.mstatus.mprv,
                         csrs.mstatus.xs,
                         csrs.mstatus.fs,
                         csrs.mstatus.mpp,
                         2b0,
                         csrs.mstatus.spp,
                         csrs.mstatus.mpie,
                         1b0,
                         csrs.mstatus.spie,
                         csrs.mstatus.upie,
                         csrs.mstatus.mie,
                         1b0,
                         csrs.mstatus.sie,
                         csrs.mstatus.uie
            );
        csr_combs.mie = bundle(20b0,
                     csrs.mie.meip,
                     1b0,
                     csrs.mie.seip,
                     csrs.mie.ueip,
                     csrs.mie.mtip,
                     1b0,
                     csrs.mie.stip,
                     csrs.mie.utip,
                     csrs.mie.msip,
                     1b0,
                     csrs.mie.ssip,
                     csrs.mie.usip );
        csr_combs.mip = bundle(20b0,
                     csrs.mip.meip,
                     1b0,
                     csrs.mip.seip,
                     csrs.mip.ueip,
                     csrs.mip.mtip,
                     1b0,
                     csrs.mip.stip,
                     csrs.mip.utip,
                     csrs.mip.msip,
                     1b0,
                     csrs.mip.ssip,
                     csrs.mip.usip );
        csr_combs.mtvec = bundle(csrs.mtvec.base, 1b0, csrs.mtvec.vectored);

        csr_combs.ustatus = bundle(27b0,
                                   csrs.mstatus.upie,
                                   3b0,
                                   csrs.mstatus.uie );
        csr_combs.uie = bundle(23b0,
                                   csrs.mie.ueip,
                                   3b0,
                                   csrs.mie.utip,
                                   3b0,
                                   csrs.mie.usip );
        csr_combs.uip = bundle(23b0,
                                   csrs.mip.ueip,
                                   3b0,
                                   csrs.mip.utip,
                                   3b0,
                                   csrs.mip.usip );
        csr_combs.utvec = bundle(csrs.utvec.base, 1b0, csrs.utvec.vectored);

        csr_combs.dcsr = bundle(csrs.dcsr.xdebug_ver,
                      12b0,
                      csrs.dcsr.ebreakm,
                      1b0,
                      csrs.dcsr.ebreaks,
                      csrs.dcsr.ebreaku,
                      csrs.dcsr.stepie,
                      csrs.dcsr.stopcount,
                      csrs.dcsr.stoptime,
                      csrs.dcsr.cause,
                      1b0,
                      csrs.dcsr.mprven,
                      csrs.dcsr.nmip,
                      csrs.dcsr.step,
                      csrs.dcsr.prv );
    }

    /*b CSR read data handling
     */
    csr_read_data """
    """: {
        /*b Decode read data */
        csr_data = {*=0};
        part_switch (csr_access.select) {
        case riscv_csr_select_time_l    : { csr_data.read_data = csrs.time[32; 0];    }
        case riscv_csr_select_time_h    : { csr_data.read_data = csrs.time[32;32];    }
        case riscv_csr_select_cycle_l   : { csr_data.read_data = csrs.cycles[32; 0];  }
        case riscv_csr_select_cycle_h   : { csr_data.read_data = csrs.cycles[32;32];  }
        case riscv_csr_select_instret_l : { csr_data.read_data = csrs.instret[32; 0]; }
        case riscv_csr_select_instret_h : { csr_data.read_data = csrs.instret[32;32]; }

        case riscv_csr_machine_isa      : { csr_data.read_data = misa      | csr_access.custom.misa;       }
        case riscv_csr_machine_vendorid : { csr_data.read_data = mvendorid | csr_access.custom.mvendorid;  }
        case riscv_csr_machine_archid   : { csr_data.read_data = marchid   | csr_access.custom.marchid;  }
        case riscv_csr_machine_impid    : { csr_data.read_data = mimpid    | csr_access.custom.mimpid;     }
        case riscv_csr_machine_hartid   : { csr_data.read_data = mhartid   | csr_access.custom.mhartid;    }

        case riscv_csr_user_status     : { csr_data.read_data = csr_combs.ustatus; }
        case riscv_csr_user_scratch    : { csr_data.read_data = csrs.uscratch; }
        case riscv_csr_user_ie         : { csr_data.read_data = csr_combs.uie; }
        case riscv_csr_user_ip         : { csr_data.read_data = csr_combs.uip; }
        case riscv_csr_user_tvec       : { csr_data.read_data = csr_combs.utvec; }
        case riscv_csr_user_tval       : { csr_data.read_data = csrs.utval; }
        case riscv_csr_user_epc        : { csr_data.read_data = csrs.uepc; }
        case riscv_csr_user_cause      : { csr_data.read_data = csrs.ucause; }

        case riscv_csr_machine_status  : { csr_data.read_data = csr_combs.mstatus; }
        case riscv_csr_machine_scratch : { csr_data.read_data = csrs.mscratch; }
        case riscv_csr_machine_ie      : { csr_data.read_data = csr_combs.mie; }
        case riscv_csr_machine_ip      : { csr_data.read_data = csr_combs.mip; }
        case riscv_csr_machine_tvec    : { csr_data.read_data = csr_combs.mtvec; }
        case riscv_csr_machine_tval    : { csr_data.read_data = csrs.mtval; }
        case riscv_csr_machine_epc     : { csr_data.read_data = csrs.mepc; }
        case riscv_csr_machine_cause   : { csr_data.read_data = csrs.mcause; }

        case riscv_csr_machine_edeleg  : { csr_data.read_data = 0; }
        case riscv_csr_machine_ideleg  : { csr_data.read_data = 0; }

        case riscv_csr_debug_pc        : { csr_data.read_data = csrs.depc; }
        case riscv_csr_debug_csr       : { csr_data.read_data = csr_combs.dcsr; }
        case riscv_csr_debug_scratch0  : { csr_data.read_data = csrs.dscratch0; }
        case riscv_csr_debug_scratch1  : { csr_data.read_data = csrs.dscratch1; }
        }
    }

    /*b CSR write controls
     */
    csr_write_controls """
    """: {
        /*b Decode CSR writes */
        csr_write.enable = 0;
        csr_write.data_mask  = 0;
        csr_write.data_set   = csr_access.write_data;
        part_switch (csr_access.access) {
            case riscv_csr_access_write: { csr_write.enable=1; }
            case riscv_csr_access_rw:    { csr_write.enable=1; }
            case riscv_csr_access_rs:    { csr_write.enable=1; csr_write.data_mask = -1; }
            case riscv_csr_access_rc:    { csr_write.enable=1; csr_write.data_set = 0; csr_write.data_mask = ~csr_access.write_data; }
        }
        if (csr_access.access_cancelled) { csr_write.enable=0; }

        /*b All done */
    }

    /*b Break out ret and trap */
    ret_trap_breakout: {
        trap_combs = {*=0};
        ret_combs = {*=0};
        if (csr_controls.trap.valid) {
            if (csr_controls.trap.ebreak_to_dbg) {
                trap_combs.d = 1;
            } elsif (csr_controls.trap.ret) {
                full_switch (csr_controls.trap.cause) {
                case riscv_trap_cause_ret_dret: { ret_combs.d = 1; }
                case riscv_trap_cause_ret_mret: { ret_combs.m = 1; }
                case riscv_trap_cause_ret_sret: { ret_combs.s = 1; }
                case riscv_trap_cause_ret_uret: { ret_combs.u = 1; }
                }
            } else {
                full_switch (csr_controls.trap.to_mode) {
                case rv_mode_debug:      { trap_combs.d = 1; }
                case rv_mode_machine:    { trap_combs.m = 1; }
                case rv_mode_supervisor: { trap_combs.s = 1; }
                case rv_mode_user:       { trap_combs.u = 1; }
                }
            }
        }
    }

    /*b CSR state update */
    csr_state_update """
    """: {
        /*b Mirror time */
        csrs.time <= irqs.time;

        /*b Handle CSR cycle state */
        csrs.cycles[32;0] <= csrs.cycles[32;0] + 1;
        if (csrs.cycles[32;0]==-1) {csrs.cycles[32;32] <= csrs.cycles[32;32]+1;}

        if (csr_write.enable && (csr_access.select==riscv_csr_select_cycle_l)) {
            csrs.cycles[32; 0]    <= (csrs.cycles[32; 0] & csr_write.data_mask) | csr_write.data_set;
        }
        if (csr_write.enable && (csr_access.select==riscv_csr_select_cycle_h)) {
            csrs.cycles[32;32]   <= (csrs.cycles[32;32] & csr_write.data_mask) | csr_write.data_set;
        }

        /*b Handle instruction retire counter state */
        if (csr_controls.retire) {
            csrs.instret[32;0] <= csrs.instret[32;0] + 1;
            if (csrs.instret[32;0]==-1) {csrs.instret[32;32] <= csrs.instret[32;32]+1;}
        }
        if (csr_write.enable && (csr_access.select==riscv_csr_select_instret_l)) {
            csrs.instret[32; 0]    <= (csrs.instret[32; 0] & csr_write.data_mask) | csr_write.data_set;
        }
        if (csr_write.enable && (csr_access.select==riscv_csr_select_instret_h)) {
            csrs.instret[32;32]   <= (csrs.instret[32;32] & csr_write.data_mask) | csr_write.data_set;
        }

        /*b Handle interrupt pending/enable state */
        csrs.mip.meip <= irqs.meip;
        csrs.mip.mtip <= irqs.mtip;
        csrs.mip.msip <= irqs.msip;
        if (csr_write.enable && (csr_access.select==riscv_csr_machine_ie)) {
            csrs.mie.meip <= (csrs.mie.meip & csr_write.data_mask[11]) | csr_write.data_set[11];
            csrs.mie.mtip <= (csrs.mie.meip & csr_write.data_mask[ 7]) | csr_write.data_set[ 7];
            csrs.mie.msip <= (csrs.mie.meip & csr_write.data_mask[ 3]) | csr_write.data_set[ 3];
        }

        /*b Handle MSTATUS.upie/uie/upp */
        if (trap_combs.u) {
            // No UPP as user mode can only trap user mode: csrs.mstatus.upp  <= 0;
            csrs.mstatus.upie <= csrs.mstatus.uie;
            csrs.mstatus.uie  <= 0;
        } else {
            if (ret_combs.u) {
                // No UPP as user mode can only trap user mode: csrs.mstatus.upp  <= 0;
                csrs.mstatus.upie <= 1;
                csrs.mstatus.uie  <= csrs.mstatus.upie;
            }
            if (csr_write.enable && (csr_access.select==riscv_csr_machine_status)) {
                // No UPP as user mode can only trap user mode: csrs.mstatus.upp <= csr_write.data[2;11];
                csrs.mstatus.upie <= (csrs.mstatus.upie & csr_write.data_mask[4]) | csr_write.data_set[4];
                csrs.mstatus.uie  <= (csrs.mstatus.uie  & csr_write.data_mask[0]) | csr_write.data_set[0];
            }
            if (csr_write.enable && (csr_access.select==riscv_csr_user_status)) {
                // No UPP as user mode can only trap user mode: csrs.mstatus.upp <= csr_write.data[2;11];
                csrs.mstatus.upie <= (csrs.mstatus.upie & csr_write.data_mask[4]) | csr_write.data_set[4];
                csrs.mstatus.uie  <= (csrs.mstatus.uie  & csr_write.data_mask[0]) | csr_write.data_set[0];
            }
        }

        /*b Handle MSTATUS.mpie/mie/mpp */
        if (trap_combs.m) {
            csrs.mstatus.mpp  <= csr_controls.exec_mode[2;0];
            csrs.mstatus.mpie <= csrs.mstatus.mie;
            csrs.mstatus.mie  <= 0;
        } else {
            if (ret_combs.m) { // note, should enter mode 'csrs.mstatus.mpp'
                csrs.mstatus.mpp  <= 0; // if machine mode only is supported, we pick that up later
                csrs.mstatus.mpie <= 1;
                csrs.mstatus.mie  <= csrs.mstatus.mpie;
            }
            if (csr_write.enable && (csr_access.select==riscv_csr_machine_status)) {
                csrs.mstatus.mpp  <= (csrs.mstatus.mpp  & csr_write.data_mask[2;11]) | csr_write.data_set[2;11];
                csrs.mstatus.mpie <= (csrs.mstatus.mpie & csr_write.data_mask[7])    | csr_write.data_set[7];
                csrs.mstatus.mie  <= (csrs.mstatus.mie  & csr_write.data_mask[3])    | csr_write.data_set[3];
            }
        }

        /*b Handle UEPC state */
        if (csr_write.enable && (csr_access.select==riscv_csr_user_epc)) {
            csrs.uepc   <= (csrs.uepc & csr_write.data_mask) | csr_write.data_set;
        }
        if (trap_combs.u) {
            csrs.uepc <= csr_controls.trap.pc;
        }

        /*b Handle MEPC state */
        if (csr_write.enable && (csr_access.select==riscv_csr_machine_epc)) {
            csrs.mepc   <= (csrs.mepc & csr_write.data_mask) | csr_write.data_set;
        }
        if (trap_combs.m) {
            csrs.mepc <= csr_controls.trap.pc;
        }

        /*b Handle DEPC state */
        if (csr_write.enable && (csr_access.select==riscv_csr_debug_pc)) {
            csrs.depc   <= (csrs.depc & csr_write.data_mask) | csr_write.data_set;
        }
        if (trap_combs.d) {
            csrs.depc <= csr_controls.trap.pc;
        }

        /*b Handle UTVEC state */
        if (csr_write.enable && (csr_access.select==riscv_csr_user_tvec)) {
            csrs.utvec.base      <= (csrs.utvec.base     & csr_write.data_mask[30;2])    | csr_write.data_set[30;2];
            csrs.utvec.vectored  <= (csrs.utvec.vectored & csr_write.data_mask[   0])    | csr_write.data_set[   0];
        }

        /*b Handle MTVEC state */
        if (csr_write.enable && (csr_access.select==riscv_csr_machine_tvec)) {
            csrs.mtvec.base      <= (csrs.mtvec.base     & csr_write.data_mask[30;2])    | csr_write.data_set[30;2];
            csrs.mtvec.vectored  <= (csrs.mtvec.vectored & csr_write.data_mask[   0])    | csr_write.data_set[   0];
        }

        /*b Handle UTVAL state */
        if (csr_write.enable && (csr_access.select==riscv_csr_user_tval)) {
            csrs.utval  <= (csrs.utval & csr_write.data_mask)    | csr_write.data_set;
        }
        if (trap_combs.u) {
            csrs.utval <= csr_controls.trap.value;
        }

        /*b Handle MTVAL state */
        if (csr_write.enable && (csr_access.select==riscv_csr_machine_tval)) {
            csrs.mtval  <= (csrs.mtval & csr_write.data_mask)    | csr_write.data_set;
        }
        if (trap_combs.m) {
            csrs.mtval <= csr_controls.trap.value;
        }

        /*b Handle UCAUSE state */
        if (csr_write.enable && (csr_access.select==riscv_csr_user_cause)) {
            csrs.ucause  <= (csrs.ucause & csr_write.data_mask)    | csr_write.data_set;
        }
        if (trap_combs.u) {
            full_switch (csr_controls.trap.cause) {
            case riscv_trap_cause_instruction_misaligned: { csrs.ucause <= bundle(24b0, riscv_mcause_instruction_misaligned); }
            case riscv_trap_cause_instruction_fault:      { csrs.ucause <= bundle(24b0, riscv_mcause_instruction_fault); }
            case riscv_trap_cause_illegal_instruction:    { csrs.ucause <= bundle(24b0, riscv_mcause_illegal_instruction); }
            case riscv_trap_cause_breakpoint:             { csrs.ucause <= bundle(24b0, riscv_mcause_breakpoint); }
            case riscv_trap_cause_load_misaligned:        { csrs.ucause <= bundle(24b0, riscv_mcause_load_misaligned); }
            case riscv_trap_cause_load_fault:             { csrs.ucause <= bundle(24b0, riscv_mcause_load_fault); }
            case riscv_trap_cause_store_misaligned:       { csrs.ucause <= bundle(24b0, riscv_mcause_store_misaligned); }
            case riscv_trap_cause_store_fault:            { csrs.ucause <= bundle(24b0, riscv_mcause_store_fault); }
            case riscv_trap_cause_uecall:                 { csrs.ucause <= bundle(24b0, riscv_mcause_uecall); }
            case riscv_trap_cause_secall:                 { csrs.ucause <= bundle(24b0, riscv_mcause_secall); }
            case riscv_trap_cause_mecall:                 { csrs.ucause <= bundle(24b0, riscv_mcause_mecall); }
            default:                                      { csrs.ucause <= bundle(1b1, 23b0, 4b0, csr_controls.trap.cause[4;0]); } // interrupts
            }
        }

        /*b Handle MCAUSE state */
        if (csr_write.enable && (csr_access.select==riscv_csr_machine_cause)) {
            csrs.mcause  <= (csrs.mcause & csr_write.data_mask)    | csr_write.data_set;
        }
        if (trap_combs.m) {
            full_switch (csr_controls.trap.cause) {
            case riscv_trap_cause_instruction_misaligned: { csrs.mcause <= bundle(24b0, riscv_mcause_instruction_misaligned); }
            case riscv_trap_cause_instruction_fault:      { csrs.mcause <= bundle(24b0, riscv_mcause_instruction_fault); }
            case riscv_trap_cause_illegal_instruction:    { csrs.mcause <= bundle(24b0, riscv_mcause_illegal_instruction); }
            case riscv_trap_cause_breakpoint:             { csrs.mcause <= bundle(24b0, riscv_mcause_breakpoint); }
            case riscv_trap_cause_load_misaligned:        { csrs.mcause <= bundle(24b0, riscv_mcause_load_misaligned); }
            case riscv_trap_cause_load_fault:             { csrs.mcause <= bundle(24b0, riscv_mcause_load_fault); }
            case riscv_trap_cause_store_misaligned:       { csrs.mcause <= bundle(24b0, riscv_mcause_store_misaligned); }
            case riscv_trap_cause_store_fault:            { csrs.mcause <= bundle(24b0, riscv_mcause_store_fault); }
            case riscv_trap_cause_uecall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_uecall); }
            case riscv_trap_cause_secall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_secall); }
            case riscv_trap_cause_mecall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_mecall); }
            default:                                      { csrs.mcause <= bundle(1b1, 23b0, 4b0, csr_controls.trap.cause[4;0]); } // interrupts
            }
        }

        /*b Handle USCRATCH state */
        if (csr_write.enable && (csr_access.select==riscv_csr_user_scratch)) {
            csrs.uscratch  <= (csrs.uscratch & csr_write.data_mask)    | csr_write.data_set;
        }

        /*b Handle MSCRATCH state */
        if (csr_write.enable && (csr_access.select==riscv_csr_machine_scratch)) {
            csrs.mscratch  <= (csrs.mscratch & csr_write.data_mask)    | csr_write.data_set;
        }

        /*b Handle DSCRATCH state */
        if (csr_write.enable && (csr_access.select==riscv_csr_debug_scratch0)) {
            csrs.dscratch0  <= (csrs.dscratch0 & csr_write.data_mask)    | csr_write.data_set;
        }
        if (csr_write.enable && (csr_access.select==riscv_csr_debug_scratch1)) {
            csrs.dscratch1  <= (csrs.dscratch1 & csr_write.data_mask)    | csr_write.data_set;
        }

        /*b Handle DCSR state */
        if (csr_write.enable && (csr_access.select==riscv_csr_debug_csr)) {
            csrs.dcsr.ebreakm   <= (csrs.dcsr.ebreakm   & csr_write.data_mask[15] ) | csr_write.data_set[15];
            csrs.dcsr.ebreaks   <= (csrs.dcsr.ebreaks   & csr_write.data_mask[13] ) | csr_write.data_set[13];
            csrs.dcsr.ebreaku   <= (csrs.dcsr.ebreaku   & csr_write.data_mask[12] ) | csr_write.data_set[12];
            csrs.dcsr.stepie    <= (csrs.dcsr.stepie    & csr_write.data_mask[11] ) | csr_write.data_set[11];
            csrs.dcsr.stopcount <= (csrs.dcsr.stopcount & csr_write.data_mask[10] ) | csr_write.data_set[10];
            csrs.dcsr.stoptime  <= (csrs.dcsr.stoptime  & csr_write.data_mask[9]  ) | csr_write.data_set[9];
            csrs.dcsr.mprven    <= (csrs.dcsr.mprven    & csr_write.data_mask[4]  ) | csr_write.data_set[4];
            csrs.dcsr.step      <= (csrs.dcsr.step      & csr_write.data_mask[2]  ) | csr_write.data_set[2];
            csrs.dcsr.prv       <= (csrs.dcsr.prv       & csr_write.data_mask[2;0]) | csr_write.data_set[2;0];
        }
        if (trap_combs.d) {
            csrs.dcsr.cause <= (csr_controls.trap.ebreak_to_dbg)?1:0; // 4=single step, 2=debugger halt
            csrs.dcsr.prv   <= csr_controls.exec_mode[2;0];
        }
        csrs.dcsr.xdebug_ver <= 4;

        /*b Kill registers if debug not enabled */
        if (rv_cfg_debug_force_disable) {
            csrs.depc <= 0;
            csrs.dscratch0 <= 0;
            csrs.dscratch1 <= 0;
            csrs.dcsr <= {*=0};
        }

        /*b Kill registers (many) if machine mode only (i.e. user mode not enabled) */
        if (!rv_cfg_user_mode_enable) {
            csrs.mstatus.mpp    <= 2b11; // only machine mode supported
            csrs.mstatus.sd     <= 0;
            csrs.mstatus.tsr    <= 0;
            csrs.mstatus.tw     <= 0;
            csrs.mstatus.tvm    <= 0;
            csrs.mstatus.mxr    <= 0;
            csrs.mstatus.sum    <= 0;
            csrs.mstatus.mprv   <= 0;
            csrs.mstatus.xs     <= 0;
            csrs.mstatus.fs     <= 0;
            csrs.mstatus.spp    <= 0;
            csrs.mstatus.spie   <= 0;
            csrs.mstatus.sie    <= 0;
            csrs.mstatus.upie   <= 0;
            csrs.mstatus.uie    <= 0;

            csrs.mip.seip     <= 0; // supervisor external interrupt pending from input pin
            csrs.mip.seip_sw  <= 0; // supervisor external interrupt pending from machine mode write
            csrs.mip.stip     <= 0; // supervisor timer interrupt pending from machine mode write
            csrs.mip.ssip     <= 0; // supervisor software interrupt pending from machine/supervisor mode write

            csrs.mie.seip     <= 0;
            csrs.mie.stip     <= 0;
            csrs.mie.ssip     <= 0;

            csrs.mip.ueip     <= 0; // user external interrupt pending from input pin
            csrs.mip.ueip_sw  <= 0; // user external interrupt pending from machine mode write
            csrs.mip.utip     <= 0; // user timer interrupt pending from machine/supervisor mode write
            csrs.mip.usip     <= 0; // user software interrupt pending from machine/supervisor mode write

            csrs.mie.ueip     <= 0;
            csrs.mie.utip     <= 0;
            csrs.mie.usip     <= 0;

            csrs.uscratch <= 0;
            csrs.uepc     <= 0;
            csrs.ucause   <= 0;
            csrs.utval    <= 0;
            csrs.utvec    <= {*=0};
        }

        /*b Kill registers (uscratch, uepc, ucause, utval, utvec) if user irq mode not enabled */
        if (!rv_cfg_user_irq_mode_enable) {
            csrs.uscratch <= 0;
            csrs.uepc     <= 0;
            csrs.ucause   <= 0;
            csrs.utval    <= 0;
            csrs.utvec    <= {*=0};
        }

        /*b Kill registers if supervisor mode not enabled */
        if (!rv_cfg_supervisor_mode_enable) {
            csrs.mstatus.spp    <= 0;
            csrs.mstatus.spie   <= 0;
            csrs.mstatus.sie    <= 0;

            csrs.mip.seip     <= 0; // supervisor external interrupt pending from input pin
            csrs.mip.seip_sw  <= 0; // supervisor external interrupt pending from machine mode write
            csrs.mip.stip     <= 0; // supervisor timer interrupt pending from machine mode write
            csrs.mip.ssip     <= 0; // supervisor software interrupt pending from machine/supervisor mode write

            csrs.mie.seip     <= 0;
            csrs.mie.stip     <= 0;
            csrs.mie.ssip     <= 0;
        }

        /*b Future - handle mtvec bounding

        The mtvec register must always be implemented, but can contain
        a hardwired read-only value. If mtvec is writable, the set of
        values the register may hold can vary by implementation. The
        value in the BASE field must always be aligned on a 4-byte
        boundary, and the MODE setting may impose additional alignment
        constraints on the value in the BASE field.

        The encoding of the MODE field is shown in Table 3.5
        (0->direct, 1->vectored, else reserved). When MODE=Direct, all
        traps into machine mode cause the pc to be set to the address
        in the BASE field. When MODE=Vectored, all synchronous
        exceptions into machine mode cause the pc to be set to the
        address in the BASE field, whereas interrupts cause the pc to
        be set to the address in the BASE field plus four times the
        interrupt cause number. For example, a machine-mode timer
        interrupt (see Table 3.6) causes the pc to be set to
        BASE+0x1c.

        Allowing coarser alignments in Vectored mode enables vectoring
        to be implemented without a hardware adder circuit.

        mtvec could be hardwired to a value - all exceptions go to
        that address (if bit 0 clear) or vectored off that address.

        Presumably utvec is similar, but should be more flexibly set
        since user mode code can occur in fewer places than machine mode.

        */

        /*b All done */
    }

    /*b Logging */
    logging """
    """: {
        if (csr_write.enable) {
            if (csr_access.address == CSR_ADDR_DSCRATCH0) {
                log("Scratch debug 0 write",
                    "write_data", csr_access.write_data );
            }
        }
    }
}


