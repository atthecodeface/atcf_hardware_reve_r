/** @copyright (C) 2016-2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 * This is a two-stage pipeline implementation, with instruction fetch
 * of the next PC occuring simultaneously with the decode, register
 * read, ALU, data read/write request, data read memory access, and
 * register update.
 *
 * The instruction memory request, then, becomes valid dependent on
 * the decode of the registered instruction last fetched. For most
 * branches this requires only a small amount of logic, but for
 * jump-and-link-register instructions (which uses the full ALU
 * result) this may take a considerable amount of gates to determine
 * the correct branch target and hence next instruction fetch.  Hence
 * the instruction memory request is valid after a considerable delay
 * from the start of the cycle.
 *
 * The return value from the instruction memory request must be valid
 * before the end of the cycle.
 *
 * Any instruction memory implementation must start its access well
 * after the CPU clock edge, , as the request is valid after the CPU
 * clock edge; the resultant read data delay (from the clock edge)
 * then has to be factored in to determine when the next CPU clock
 * edge can occur. Hence it may be sensible to use a double speed
 * clock (e.g. 'fast_clk') to generate CPU clock edges (every other
 * fast_clk edge) and SRAM access clock edges (for a synchronous
 * memory) on the intervening fast_clk edges.
 *
 * The data memory request becomes valid, again, a fair time after the
 * CPU clock edge, as it requires instruction decode, register fetch,
 * and ALU operation to occur prior to the memory address being valid.
 *
 * The data memory response must be valid (for read data!) in the same
 * CPU cycle, as the returning data has to be rotated to the correct
 * byte lanes and prepared for the register file write.
 *
 * Hence a data memory implementation can be similar to that proposed
 * for the instruction memory - that is, accesses start on a memory
 * clock edge that is in the middle of a CPU clock edge, by using a
 * fast_clk.
 *
 */

/*a Includes
 */
include "reve_r.h"
include "reve_r_fetch.h"           // for fetch request
include "reve_r_pipeline_types.h"  // for pipeline control, response, fetch_data

/*a Constants
 */
constant integer INITIAL_PC=0x0;
constant integer i32_enable_branch_prediction=1;

/*a Types
 */
/*t t_ifetch_combs
 *
 * Combinatorials for the instruction fetch
 */
typedef struct {
    bit[32] pc_plus_4;
    bit[32] pc_plus_2;
    bit[32] pc_plus_inst;
    bit[32] pc_if_mispredicted;
    bit predict_branch;
    bit[32] fetch_next_pc;
    bit     fetch_sequential;
} t_ifetch_combs;

/*a Module
 */
module reve_r_pipeline_control_fetch_req( input t_reve_r_pipeline_state        pipeline_state,
                                             input t_reve_r_pipeline_response     pipeline_response,
                                             output t_reve_r_pipeline_fetch_req   pipeline_fetch_req,
                                             output t_reve_r_fetch_req            ifetch_req
)
{
    comb t_ifetch_combs ifetch_combs;

    /*b Pipeline control
     */
    pipeline_state_logic
    """
    The instruction fetch request derives from the
    decode/execute stage (the instruction address that is required
    next) and presents that to the outside world.

    This request may be for any 16-bit aligned address, and two
    successive 16-bit words from that request must be presented,
    aligned to bit 0.

    If the decode/execute stage is invalid (i.e. it does not have a
    valid instruction to decode) then the current PC is requested.
    """:
    {
        //ifetch_combs.pc_plus_4     = pipeline_state.fetch_pc + 4;
        //ifetch_combs.pc_plus_2     = pipeline_state.fetch_pc + 2;
        ifetch_combs.pc_plus_4     = pipeline_response.decode.pc + 4;
        ifetch_combs.pc_plus_2     = pipeline_response.decode.pc + 2;
        ifetch_combs.pc_plus_inst  = ifetch_combs.pc_plus_4;
        if (pipeline_response.decode.idecode.is_compressed) {
            ifetch_combs.pc_plus_inst = ifetch_combs.pc_plus_2;
        }

        /*b Detect unconditional branches and backward conditional branches */
        ifetch_combs.predict_branch    = 0;
        part_switch (pipeline_response.decode.idecode.op) {
        case reve_r_op_branch:   { ifetch_combs.predict_branch = pipeline_response.decode.idecode.immediate[31]; }
        case reve_r_op_jal:      { ifetch_combs.predict_branch = 1; }
        }
        if (rv_cfg_i32c_force_disable /*|| !riscv_config.i32c */) {
            if (pipeline_response.decode.branch_target[1]) {
                ifetch_combs.predict_branch = 0;
            }
        }
        if (!i32_enable_branch_prediction || !pipeline_response.decode.enable_branch_prediction) {
            ifetch_combs.predict_branch = 0;
        }

        ifetch_combs.fetch_next_pc      = ifetch_combs.pc_plus_inst;
        ifetch_combs.fetch_sequential   = 1;
        ifetch_combs.pc_if_mispredicted = pipeline_response.decode.branch_target;
        if (ifetch_combs.predict_branch) {
            ifetch_combs.fetch_next_pc      = pipeline_response.decode.branch_target;
            ifetch_combs.fetch_sequential   = 0;
            ifetch_combs.pc_if_mispredicted = ifetch_combs.pc_plus_inst;
        }

        /*b Determine ifetch_req and pipeline_fetch_req */
        ifetch_req                 = {*=0};
        pipeline_fetch_req         = {*=0};

        pipeline_fetch_req.predicted_branch   = ifetch_combs.predict_branch;
        pipeline_fetch_req.pc_if_mispredicted = ifetch_combs.pc_if_mispredicted;
        ifetch_req.flush_pipeline = 1;
        ifetch_req.req_type = rv_fetch_none;
        ifetch_req.address  = pipeline_state.fetch_pc; // == ifetch_state.pc
        ifetch_req.mode     = pipeline_state.mode;

        full_switch (pipeline_state.fetch_action) {
        case rv_pc_fetch_action_restart_at_pc: {
            ifetch_req.flush_pipeline = 1;
            ifetch_req.req_type       = rv_fetch_nonsequential;
            ifetch_req.address        = pipeline_state.fetch_pc;
        }
        case rv_pc_fetch_action_retry: {
            ifetch_req.flush_pipeline = 0;
            ifetch_req.req_type       = rv_fetch_repeat;
            ifetch_req.address        = pipeline_state.fetch_pc;
        }
        case rv_pc_fetch_action_continue_fetching: {
            ifetch_req.flush_pipeline = 0;
            ifetch_req.req_type       = rv_fetch_nonsequential;
            if (ifetch_combs.fetch_sequential) {
                ifetch_req.req_type = (pipeline_response.decode.idecode.is_compressed) ? rv_fetch_sequential_16 : rv_fetch_sequential_32;
            }
            ifetch_req.address        = ifetch_combs.fetch_next_pc; // early address
        }
        case rv_pc_fetch_action_none: {
            ifetch_req.flush_pipeline = 0;
        }
        default: { // idle
            ifetch_req.flush_pipeline = 1;
        }
        }

        pipeline_fetch_req.debug_fetch = 0;
        if (pipeline_state.mode == rv_mode_debug) {
            if ((pipeline_state.fetch_action!=rv_pc_fetch_action_idle) &&
                (pipeline_state.fetch_action!=rv_pc_fetch_action_none) &&
                (ifetch_req.address[24;8]==-1)) {
                ifetch_req.req_type = rv_fetch_none;
                ifetch_req.mode     = rv_mode_debug;
                pipeline_fetch_req.debug_fetch = 1;
            }
        }

        /*b All done
         */
    }
}
