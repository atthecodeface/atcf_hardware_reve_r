/** @copyright (C) 2018-2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_pipeline_debug.cdl
 * @brief  Low-gate-count RISC-V pipeline debug module
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 */

/*a Includes
 */
include "reve_r.h"
include "reve_r_fetch.h"           // for fetch request
include "reve_r_pipeline_types.h"  // for pipeline debug control, response
include "reve_r_debug.h"

/*a Constants
 */

/*a Types
 */
/*t t_debug_fsm
 *
 * State machine
 */
typedef fsm {
    debug_fsm_running;
    debug_fsm_halting;
    debug_fsm_halted;
    debug_fsm_resuming;
        
    // runnning, halting, resuming, single step, read register_start, read_register_wait, write register_start, write_register_wait, 
} t_debug_fsm;

/*t t_debug_combs
 *
 * Combinatorial signals from the state and inputs
 *
 */
typedef struct {
    bit mst_valid;
} t_debug_combs;

/*t t_debug_state
 *
 * State of debugger 
 *
 */
typedef struct {
    t_debug_fsm fsm_state;
    bit drive_attention;
    bit drive_response;
    bit halt_req;
    bit resume_req;
    bit halted;
    bit resumed;
    bit attention;
    bit hit_breakpoint;
    bit[16] arg;
    bit[6] rv_select;
    t_reve_r_debug_resp resp "Response from a requested op - only one op should be requested for each response";
    bit[32] data0      "Data from a completed transaction; 0 otherwise";
} t_debug_state;

/*a Module
 */
module reve_r__pipeline_debug( clock clk,
                                 input bit reset_n,
                                 input  t_reve_r_debug_mst debug_mst,
                                 output t_reve_r_debug_tgt debug_tgt,
                                 output t_reve_r_pipeline_debug_control debug_control,
                                 input  t_reve_r_pipeline_debug_response debug_response,

                                 input bit[6] rv_select
)
"""
This is a fully synchronous pipeline debug module. 

It is designed to feed data in to a RISC-V pipeline (being merged with
instruction fetch responses), and it takes commands and reports out to
a RISC-V debug module.

"""
{

    /*b State and comb
     */
    default clock clk;
    default reset active_low reset_n;

    comb t_debug_combs debug_combs;
    clocked t_debug_state debug_state = {*=0};

    /*b Drive control of the pipeline
     */
    pipeline_control """
    """ : {
        debug_control = {*=0};
        debug_control.valid = 0;
        debug_control.data  = debug_state.data0;
        debug_control.kill_fetch = 0;
        debug_control.halt_request = 0; // forces entry to debug mode
        full_switch (debug_state.fsm_state) {
        case debug_fsm_running: {
            debug_control.kill_fetch = 0;
        }
        case debug_fsm_halting: {
            debug_control.valid = 1;
            debug_control.kill_fetch = 1;
            debug_control.halt_request = 1; // forces entry to debug mode
        }
        case debug_fsm_halted: {
            debug_control.valid = 1;
            debug_control.kill_fetch = 1;
        }
        case debug_fsm_resuming: {
            debug_control.valid = 1;
            debug_control.fetch_dret = 1; // forces a dret?
        }
        }
    }

    /*b Debug state machine
     */
    debug_state_machine """
    """ : {
        debug_combs.mst_valid = debug_mst.valid;
        if (debug_mst.select != rv_select) {
            debug_combs.mst_valid = 0;
        }
        if (debug_combs.mst_valid) {
            debug_state.attention <= 0;
            if (debug_mst.op==rv_debug_set_requests) {
                debug_state.halt_req <= debug_mst.arg[0];
                debug_state.resume_req <= debug_mst.arg[1];
            }
            if (debug_mst.op==rv_debug_read) {
                debug_state.arg   <= debug_mst.arg;
                debug_state.data0 <= debug_mst.data;
            }
        }

        debug_state.resp <= {*=0};
        if (debug_state.resumed && !debug_state.resume_req) {
            debug_state.resumed <= 0;
            debug_state.attention <= 1;
        }

        full_switch (debug_state.fsm_state) {
        case debug_fsm_running: {
            if (debug_state.halt_req) {
                debug_state.fsm_state <= debug_fsm_halting;
            }
            if (debug_response.exec_valid && debug_response.exec_halting) { // ebreak?
                debug_state.fsm_state <= debug_fsm_halted;
                debug_state.halted <= 1;
                debug_state.hit_breakpoint <= 1;
                debug_state.attention <= 1;
            }
        }
        case debug_fsm_halting: {
            if (debug_response.exec_valid && debug_response.exec_halting) {
                debug_state.fsm_state <= debug_fsm_halted;
                debug_state.halted <= 1;
                debug_state.attention <= 1;
            }
        }
        case debug_fsm_halted: { // can resume or single step from here (or read/write register, or execute progbuf)
            if (debug_state.resume_req && !debug_state.resumed) {
                debug_state.fsm_state <= debug_fsm_resuming;
            }
        }
        case debug_fsm_resuming: {
            if (debug_response.exec_valid && debug_response.exec_dret) {
                debug_state.fsm_state <= debug_fsm_running;
                debug_state.hit_breakpoint <= 0;
                debug_state.halted <= 0;
                debug_state.resumed <= 1;
                debug_state.attention <= 1;
            }
        }
        }
    }

    /*b Drive debug response
     */
    debug_response_driving """
    """ : {

        debug_state.drive_attention <= 0;
        debug_state.drive_response  <= 0;
        if ((debug_mst.mask & rv_select) == debug_mst.select) {
            debug_state.drive_attention <= 1;
        }
        if (debug_mst.valid && (rv_select==debug_mst.select)) {
            debug_state.drive_response <= 1;
        }
        if (debug_state.rv_select!=0) {
            debug_state.rv_select <= rv_select;
        }

        debug_tgt = {*=0};
        if (debug_state.drive_attention) {
            debug_tgt.attention = debug_state.attention;
        }
        if (debug_state.drive_response) {
            debug_tgt.valid          = 1;
            debug_tgt.selected       = debug_state.rv_select;
            debug_tgt.halted         = debug_state.halted;
            debug_tgt.resumed        = debug_state.resumed;
            debug_tgt.hit_breakpoint = debug_state.hit_breakpoint;
            debug_tgt.resp           = debug_state.resp;
            debug_tgt.data           = debug_state.data0;
        }
    }
}
