/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 * This is a two-stage pipeline implementation, with instruction fetch
 * of the next PC occuring simultaneously with the decode, register
 * read, ALU, data read/write request, data read memory access, and
 * register update.
 *
 * The instruction memory request, then, becomes valid dependent on
 * the decode of the registered instruction last fetched. For most
 * branches this requires only a small amount of logic, but for
 * jump-and-link-register instructions (which uses the full ALU
 * result) this may take a considerable amount of gates to determine
 * the correct branch target and hence next instruction fetch.  Hence
 * the instruction memory request is valid after a considerable delay
 * from the start of the cycle.
 *
 * The return value from the instruction memory request must be valid
 * before the end of the cycle.
 *
 * Any instruction memory implementation must start its access well
 * after the CPU clock edge, , as the request is valid after the CPU
 * clock edge; the resultant read data delay (from the clock edge)
 * then has to be factored in to determine when the next CPU clock
 * edge can occur. Hence it may be sensible to use a double speed
 * clock (e.g. 'fast_clk') to generate CPU clock edges (every other
 * fast_clk edge) and SRAM access clock edges (for a synchronous
 * memory) on the intervening fast_clk edges.
 *
 * The data memory request becomes valid, again, a fair time after the
 * CPU clock edge, as it requires instruction decode, register fetch,
 * and ALU operation to occur prior to the memory address being valid.
 *
 * The data memory response must be valid (for read data!) in the same
 * CPU cycle, as the returning data has to be rotated to the correct
 * byte lanes and prepared for the register file write.
 *
 * Hence a data memory implementation can be similar to that proposed
 * for the instruction memory - that is, accesses start on a memory
 * clock edge that is in the middle of a CPU clock edge, by using a
 * fast_clk.
 *
 */

/*a Includes
 */
include "reve_r.h"
include "reve_r_fetch.h"           // for fetch request
include "reve_r_pipeline_types.h"  // for pipeline control, response, fetch_data

/*a Module
 */
module reve_r_pipeline_control_fetch_data( input t_reve_r_pipeline_state       pipeline_state,
                                              input  t_reve_r_fetch_req           ifetch_req,
                                              input  t_reve_r_fetch_resp          ifetch_resp,
                                              input t_reve_r_pipeline_fetch_req   pipeline_fetch_req,
                                              output t_reve_r_pipeline_fetch_data pipeline_fetch_data
)
{
    /*b Pipeline control
     */
    pipeline_state_logic
    """
    The instruction fetch request derives from the
    decode/execute stage (the instruction address that is required
    next) and presents that to the outside world.

    This request may be for any 16-bit aligned address, and two
    successive 16-bit words from that request must be presented,
    aligned to bit 0.

    If the decode/execute stage is invalid (i.e. it does not have a
    valid instruction to decode) then the current PC is requested.
    """:
    {
        pipeline_fetch_data.valid = ifetch_resp.valid && (ifetch_req.req_type != rv_fetch_none);
        pipeline_fetch_data.pc    = ifetch_req.address;
        pipeline_fetch_data.mode  = ifetch_req.mode;
        pipeline_fetch_data.instruction  = {data=ifetch_resp.data, mode=ifetch_req.mode, debug={*=0}};
        if (pipeline_fetch_req.debug_fetch) {
            if (ifetch_req.address[8;0]==0) {
                pipeline_fetch_data.valid = 1;
                pipeline_fetch_data.instruction.data=pipeline_state.instruction_data;
            } else {
                pipeline_fetch_data.valid = 1;
                pipeline_fetch_data.instruction.data=RV32I_EBREAK;
            }
        }
        pipeline_fetch_data.dec_pc_if_mispredicted = pipeline_fetch_req.pc_if_mispredicted;
        pipeline_fetch_data.dec_predicted_branch   = pipeline_fetch_req.predicted_branch;

        if (pipeline_state.instruction_debug.valid) {
            pipeline_fetch_data.valid = 1;
            pipeline_fetch_data.instruction.debug  = pipeline_state.instruction_debug;
            pipeline_fetch_data.instruction.data   = pipeline_state.instruction_data;
        }
    }
}
